`timescale 1ns/100ps

module immediateGenerator (
    input [32:0] instruction,
    output [11:0] immediate
);

    
endmodule