module riscv (
    input wire semente,
    input wire clock
);

    
endmodule