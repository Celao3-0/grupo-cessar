module xor (
    input [31:0] A,
    input [31:0] B,
    output [31:0] result
);
    xor (result, A, B);
endmodule