module or (
    input [31:0] A,
    input [31:0] B,
    output [31:0] result
);
    or (result, A, B);
endmodule