module riscv (
    input wire semente,
    input wire clk
);

    
endmodule