module and (
    input [31:0] A,
    input [31:0] B,
    output [31:0] result
);
    and (result, A, B);
endmodule